    module mux4(i0,i1,i2,i3,sel,out);
    input [-1:0] i0;
    input [-1:0] i1;
    input [-1:0] i2;
    input [-1:0] i3;
    input [1:0] sel;
    output [-1:0] out;
    
    assign out = ;

    endmodule
