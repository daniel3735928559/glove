    module imm_prep(c_imm_type,inst_in,imm);
    input [2:0] c_imm_type;
    input [15:0] inst_in;
    output [7:0] imm;
    
    assign imm = ;

    endmodule
