    module alu(A,B,op,T,C,result,flags);
    input [7:0] A;
    input [7:0] B;
    input [3:0] op;
    input T;
    input C;
    output [7:0] result;
    output [6:0] flags;
    
    assign result = ;
    assign flags = ;

    endmodule
