    module control(inst,state,c_new_sreg_sel,c_imem_addr_sel,c_adiw_phase,c_sp_op,c_ram_adr_sel,c_io_op,c_ram_op,c_rd_w_en,c_dbus_addr_sel,c_pc_offset_mode,c_flags_mask,c_imm_type,c_alu_b_sel,c_pc_stall,c_alu_op,c_rh_sel,c_rampz_inc,c_ex_out_sel,c_pc_next,c_rh_op,c_dbus_out_sel,c_alu_a_sel,c_mem_out_sel,c_branch_mode,c_rd_rr_sel,c_next_state,c_skip);
    input [15:0] inst;
    input [1:0] state;
    output c_new_sreg_sel;
    output [1:0] c_imem_addr_sel;
    output c_adiw_phase;
    output [1:0] c_sp_op;
    output [2:0] c_ram_adr_sel;
    output [1:0] c_io_op;
    output [1:0] c_ram_op;
    output c_rd_w_en;
    output [1:0] c_dbus_addr_sel;
    output c_pc_offset_mode;
    output [7:0] c_flags_mask;
    output [2:0] c_imm_type;
    output c_alu_b_sel;
    output c_pc_stall;
    output [3:0] c_alu_op;
    output [1:0] c_rh_sel;
    output c_rampz_inc;
    output c_ex_out_sel;
    output [2:0] c_pc_next;
    output [1:0] c_rh_op;
    output [1:0] c_dbus_out_sel;
    output [1:0] c_alu_a_sel;
    output c_mem_out_sel;
    output c_branch_mode;
    output [1:0] c_rd_rr_sel;
    output [1:0] c_next_state;
    output c_skip;
    
    assign c_new_sreg_sel = ;
    assign c_imem_addr_sel = ;
    assign c_adiw_phase = ;
    assign c_sp_op = ;
    assign c_ram_adr_sel = ;
    assign c_io_op = ;
    assign c_ram_op = ;
    assign c_rd_w_en = ;
    assign c_dbus_addr_sel = ;
    assign c_pc_offset_mode = ;
    assign c_flags_mask = ;
    assign c_imm_type = ;
    assign c_alu_b_sel = ;
    assign c_pc_stall = ;
    assign c_alu_op = ;
    assign c_rh_sel = ;
    assign c_rampz_inc = ;
    assign c_ex_out_sel = ;
    assign c_pc_next = ;
    assign c_rh_op = ;
    assign c_dbus_out_sel = ;
    assign c_alu_a_sel = ;
    assign c_mem_out_sel = ;
    assign c_branch_mode = ;
    assign c_rd_rr_sel = ;
    assign c_next_state = ;
    assign c_skip = ;

    endmodule
