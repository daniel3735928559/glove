    module inc(input,output);
    input [-1:0] input;
    output [-1:0] output;
    
    assign output = ;

    endmodule
