    module register(d,clk,rst,q);
    input [-1:0] d;
    input clk;
    input rst;
    output [-1:0] q;
    
    assign q = ;

    endmodule
