    module is_zero(d,result);
    input [-1:0] d;
    output result;
    
    assign result = (d==0);

    endmodule
