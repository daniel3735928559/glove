    module bitwise_mux(i0,i1,mask,output);
    input [7:0] i0;
    input [7:0] i1;
    input [7:0] mask;
    output [7:0] output;
    
    assign output = ;

    endmodule
