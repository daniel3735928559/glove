    module z_adder(i0,i1,output);
    input [15:0] i0;
    input [7:0] i1;
    output [15:0] output;
    
    assign output = ;

    endmodule
