    module offset_comp(pc,inst,c_pc_offset_mode,pc_plus_offset);
    input [15:0] pc;
    input [15:0] inst;
    input c_pc_offset_mode;
    output [15:0] pc_plus_offset;
    
    assign pc_plus_offset = ;

    endmodule
