    module mux2(i0,i1,sel,out);
    input [-1:0] i0;
    input [-1:0] i1;
    input sel;
    output [-1:0] out;
    
    assign out = ;

    endmodule
