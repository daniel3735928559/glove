    module is_32_bit(inst_in,is_32_bit);
    input [15:0] inst_in;
    output is_32_bit;
    
    assign is_32_bit = ;

    endmodule
