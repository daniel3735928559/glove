    module mux8(i0,i1,i2,i3,i4,i5,i6,i7,sel,out);
    input [-1:0] i0;
    input [-1:0] i1;
    input [-1:0] i2;
    input [-1:0] i3;
    input [-1:0] i4;
    input [-1:0] i5;
    input [-1:0] i6;
    input [-1:0] i7;
    input [2:0] sel;
    output [-1:0] out;
    
    assign out = ;

    endmodule
  
