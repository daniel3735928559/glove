    module loc_io_reg_file(c_rampz0_inc,dbusin,dbus_adr,sreg_in,dbus_out,sp_op,io_op,clk,rst,sreg,spl,sph,rampz,dbusin_int);
    input c_rampz0_inc;
    input [7:0] dbusin;
    input [5:0] dbus_adr;
    input [7:0] sreg_in;
    input [7:0] dbus_out;
    input [1:0] sp_op;
    input [1:0] io_op;
    input clk;
    input rst;
    output [7:0] sreg;
    output [7:0] spl;
    output [7:0] sph;
    output rampz;
    output [7:0] dbusin_int;
    
    assign sreg = ;
    assign spl = ;
    assign sph = ;
    assign rampz = ;
    assign dbusin_int = ;

    endmodule
